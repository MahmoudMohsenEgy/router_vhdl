grayCounterTestBench.vhdl
